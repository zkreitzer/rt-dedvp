// This is an example/template file in fpga/src/.
// Files in this directory implement FPGA HDL modules for the ASOC interface,
// data acquisition, buffering, and control logic.
// Replace this file with real design modules or copy/rename it when creating
// new top-level or leaf modules.

module asoc_fpga_top_example (
    input  wire clk,
    input  wire rst_n
    // TODO: add ASOC, MCP, and I/O ports
);
    // TODO: implement ASOC interface and readout logic.
endmodule

